<dec f='halide/build/_deps/pybind11-src/include/pybind11/cast.h' l='214' type='void **'/>
<use f='halide/build/_deps/pybind11-src/include/pybind11/cast.h' l='219' u='w' c='_ZN8pybind116detail16value_and_holderC1EPNS0_8instanceEPKNS0_9type_infoEmm'/>
<use f='halide/build/_deps/pybind11-src/include/pybind11/cast.h' l='229' u='r' c='_ZNK8pybind116detail16value_and_holder9value_ptrEv'/>
<use f='halide/build/_deps/pybind11-src/include/pybind11/cast.h' l='235' u='r' c='_ZNK8pybind116detail16value_and_holder6holderEv'/>
<use f='halide/build/_deps/pybind11-src/include/pybind11/cast.h' l='295' u='w' c='_ZN8pybind116detail18values_and_holders8iteratorppEv'/>
<offset>192</offset>
